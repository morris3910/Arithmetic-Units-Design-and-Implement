module HA(
    input a, b, 
    output s, c
);
  assign s = a ^ b;
  assign c = a & b;
endmodule

module FA(
    input a, b, cin, 
    output s, c
);
  assign s = a ^ b ^ cin;
  assign c = (a & b) | (b & cin) | (a & cin);
endmodule

module array_mul_8x8 (
    input [7:0] a,
    input [7:0] b,
    output [15:0] p
);
    wire [64:0] s, c;
    assign p[0] = a[0] & b[0];

    HA ha11 ((a[0] & b[1]), (a[1] & b[0]), p[1], c[0]);
    FA fa11 ((a[1] & b[1]), (a[2] & b[0]), c[0], s[1], c[1]);
    FA fa12 ((a[2] & b[1]), (a[3] & b[0]), c[1], s[2], c[2]);
    FA fa13 ((a[3] & b[1]), (a[4] & b[0]), c[2], s[3], c[3]);
    FA fa14 ((a[4] & b[1]), (a[5] & b[0]), c[3], s[4], c[4]);
    FA fa15 ((a[5] & b[1]), (a[6] & b[0]), c[4], s[5], c[5]);
    FA fa16 ((a[6] & b[1]), (a[7] & b[0]), c[5], s[6], c[6]);
    HA ha12 (c[6], (a[7] & b[1]), s[7], c[7]);

    HA ha21 ((a[0] & b[2]), s[1], p[2], c[8]);
    FA fa21 ((a[1] & b[2]), s[2], c[8], s[9], c[9]);
    FA fa22 ((a[2] & b[2]), s[3], c[9], s[10], c[10]);
    FA fa23 ((a[3] & b[2]), s[4], c[10], s[11], c[11]);
    FA fa24 ((a[4] & b[2]), s[5], c[11], s[12], c[12]);
    FA fa25 ((a[5] & b[2]), s[6], c[12], s[13], c[13]);
    FA fa26 ((a[6] & b[2]), s[7], c[13], s[14], c[14]);
    FA fa27 ((a[7] & b[2]), c[7], c[14], s[15], c[15]);

    HA ha31 ((a[0] & b[3]), s[9], p[3], c[16]);
    FA fa31 ((a[1] & b[3]), s[10], c[16], s[17], c[17]);
    FA fa32 ((a[2] & b[3]), s[11], c[17], s[18], c[18]);
    FA fa33 ((a[3] & b[3]), s[12], c[18], s[19], c[19]);
    FA fa34 ((a[4] & b[3]), s[13], c[19], s[20], c[20]);
    FA fa35 ((a[5] & b[3]), s[14], c[20], s[21], c[21]);
    FA fa36 ((a[6] & b[3]), s[15], c[21], s[22], c[22]);
    FA fa37 ((a[7] & b[3]), c[15], c[22], s[23], c[23]);

    HA ha41 ((a[0] & b[4]), s[17], p[4], c[24]);
    FA fa41 ((a[1] & b[4]), s[18], c[24], s[25], c[25]);
    FA fa42 ((a[2] & b[4]), s[19], c[25], s[26], c[26]);
    FA fa43 ((a[3] & b[4]), s[20], c[26], s[27], c[27]);
    FA fa44 ((a[4] & b[4]), s[21], c[27], s[28], c[28]);
    FA fa45 ((a[5] & b[4]), s[22], c[28], s[29], c[29]);
    FA fa46 ((a[6] & b[4]), s[23], c[29], s[30], c[30]);
    FA fa47 ((a[7] & b[4]), c[23], c[30], s[31], c[31]);

    HA ha51 ((a[0] & b[5]), s[25], p[5], c[32]);
    FA fa51 ((a[1] & b[5]), s[26], c[32], s[33], c[33]);
    FA fa52 ((a[2] & b[5]), s[27], c[33], s[34], c[34]);
    FA fa53 ((a[3] & b[5]), s[28], c[34], s[35], c[35]);
    FA fa54 ((a[4] & b[5]), s[29], c[35], s[36], c[36]);
    FA fa55 ((a[5] & b[5]), s[30], c[36], s[37], c[37]);
    FA fa56 ((a[6] & b[5]), s[31], c[37], s[38], c[38]);
    FA fa57 ((a[7] & b[5]), c[31], c[38], s[39], c[39]);

    HA ha61 ((a[0] & b[6]), s[33], p[6], c[40]);
    FA fa61 ((a[1] & b[6]), s[34], c[40], s[41], c[41]);
    FA fa62 ((a[2] & b[6]), s[35], c[41], s[42], c[42]);
    FA fa63 ((a[3] & b[6]), s[36], c[42], s[43], c[43]);
    FA fa64 ((a[4] & b[6]), s[37], c[43], s[44], c[44]);
    FA fa65 ((a[5] & b[6]), s[38], c[44], s[45], c[45]);
    FA fa66 ((a[6] & b[6]), s[39], c[45], s[46], c[46]);
    FA fa67 ((a[7] & b[6]), c[39], c[46], s[47], c[47]);

    HA ha71 ((a[0] & b[7]), s[41], p[7], c[48]);
    FA fa71 ((a[1] & b[7]), s[42], c[48], p[8], c[49]);
    FA fa72 ((a[2] & b[7]), s[43], c[49], p[9], c[50]);
    FA fa73 ((a[3] & b[7]), s[44], c[50], p[10], c[51]);
    FA fa74 ((a[4] & b[7]), s[45], c[51], p[11], c[52]);
    FA fa75 ((a[5] & b[7]), s[46], c[52], p[12], c[53]);
    FA fa76 ((a[6] & b[7]), s[47], c[53], p[13], c[54]);
    FA fa77 ((a[7] & b[7]), c[47], c[54], p[14], p[15]);

endmodule

